

library IEEE;
use IEEE.STD_LOGIC_1164.ALL; 

entity control_logic_tb is 

    
end control_logic_tb ;